`ifndef _inst
`define _inst

`define NOP 0
`define ADD 1
`define SUB 2
`define AND 3
`define OR 4
`define XOR 5

module I();endmodule

`endif
